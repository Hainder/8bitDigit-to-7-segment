module AsciiToSevenSeg (
	input [7:0] ascii,
	output [7:0] sevenSeg
);



endmodule 